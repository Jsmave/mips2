module ID_EX (
    ports
);
    
endmodule