`include "../define.v"
module EX_MEM (
    ports
);
    
endmodule