module MEM_WR (
    ports
);
    
endmodule