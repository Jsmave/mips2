`include "../define.v"
module MEM_WR (
    ports
);
    
endmodule