module mips_top_sim (

);
    
endmodule