`include "define.v"
module ControlUnit (
    input [`N:0] instruction_D,
    output wire [4:0] AluOP,
    output wire [`N:0] ControlSignal
);
    wire reg_we,ram_we;
    
    assign 
endmodule