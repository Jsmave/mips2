`include "../define.v"
module EX_MEM (
    
);
    
endmodule